module table_test
