module store_register(input wire [20:0] in, input wire [20:0] mem [20:0]);


